struct HelloWorld
{
	string msg;
};
struct PostData
{
	long a;
	long b;
};

port MyData PostData;
port OriginalData HelloWorld;
interface ADD
{
	double add(inout HelloWorld a);
};
interface MINUS
{
	double minus(in double a,out double b);
};

service component Transformer
{
	publish OriginalData OriginData1;
	provide ADD PolarUnit1;
	provide MINUS PolarUnit3;
};
ui component Sensor
{
	publish MyData TestData1;
	consume OriginalData OriginData2;
	require ADD PolarUnit2;
};
ui component Navidisplay
{
	consume MyData TestData2;
	require MINUS PolarUnit4;
};
